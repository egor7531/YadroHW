//----------------------------------------------------------------------------
// Task
//----------------------------------------------------------------------------

module round_robin_arbiter_with_2_requests
(
    input        clk,
    input        rst,
    input  [1:0] requests,
    output [1:0] grants
);

    logic [1:0] ng;
    logic[1:0] g;

    always_ff @(posedge clk) begin
        if(rst) begin
            ng <= 2'b00;
        end else begin
            ng <= requests;
        end
    end

    always_comb begin
        if(requests == 2'b11) begin
            if(~ng[0])
            g = 2'b01;
            else
            g = 2'b10;
        end else begin
            g = requests;
        end
    end

    assign grants = g;
    // Task:
    // Implement a "arbiter" module that accepts up to two requests
    // and grants one of them to operate in a round-robin manner.
    //
    // The module should maintain an internal register
    // to keep track of which requester is next in line for a grant.
    //
    // Note:
    // Check the waveform diagram in the README for better understanding.
    //
    // Example:
    // requests -> 01 00 10 11 11 00 11 00 11 11
    // grants   -> 01 00 10 01 10 00 01 00 10 01


endmodule
